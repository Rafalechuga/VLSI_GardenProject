LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--selSs7 ss70, ss71, sel, ss7Out
ENTITY selSs7 IS
PORT(
	ss70, ss71: STD_LOGIC_VECTOR( 6 DOWNTO 0 );
	sel: INTEGER RANGE 0 TO 3;
	ss7Out: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0 )
);
END ENTITY;

ARCHITECTURE arq OF selSs7 IS
BEGIN 
	WITH sel SELECT ss7Out <=
	ss70 WHEN 0,
	ss70 WHEN 1,
	ss70 WHEN 2,
	ss71 WHEN 3,
	ss71 WHEN OTHERS;		
END ARCHITECTURE;